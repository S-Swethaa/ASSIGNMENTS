`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/27/2025 09:44:46 PM
// Design Name: 
// Module Name: question_15
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module question_15();
reg [3:0]a= 4'b110x;
initial
begin
if ( a !== 4'b1100)
begin: B1
end
else
begin: B2 end
end

endmodule
