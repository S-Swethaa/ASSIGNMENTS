`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module TASK_FN_qn7_tb;
reg [4:0]x;
wire[4:0]y;
TASK_FN_qn7 u1(.y(y),.x(x));
initial begin
x=5'b11011;#10;
$finish;
end
endmodule
